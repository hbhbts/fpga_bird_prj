//utils_pkg
`ifndef UTILS_PKG_SV
`define UTILS_PKG_SV
package utils_pkg;
	parameter VERSION = 0;
endpackage
`endif

import utils_pkg::*;





