//utils_pkg
`ifndef UTILS_PKG_SV
`define UTILS_PKG_SV
package utils_pkg;
	parameter VERSION = "1.0";
endpackage

import utils_pkg::*;

`endif




